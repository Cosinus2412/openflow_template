/**
 * Package: cipher_pkg
 *
 * Defines parameters, types and conversion functions for your cipher.
 *
 */

package cipher_pkg;
  // --------------------------------------------------------------------------
  // Type definitions
  // --------------------------------------------------------------------------

  // Length definitions for the cipher
  parameter KEY_LENGTH  = 128;
  parameter DATA_LENGTH = 128;
  parameter LENGTH      = 32;
endpackage
